module CPU_Demo(
    input src_clk,
    output	[6:0] HEX0,
    output	[6:0] HEX1,
    output	[6:0] HEX2,
    output	[6:0] HEX3,
    output	[6:0] HEX4,
    output	[6:0] HEX5,
    output	[6:0] HEX6,	
    output	[6:0] HEX7 
);

reg [31:0] disp=32'h00c00193;

Digits digits(
    .disp(disp),
    
    .HEX0(HEX0),
    .HEX1(HEX1),
    .HEX2(HEX2),
    .HEX3(HEX3),

    .HEX4(HEX4),
    .HEX5(HEX5),
    .HEX6(HEX6),
    .HEX7(HEX7)
);

endmodule