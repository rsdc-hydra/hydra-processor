`ifndef PARAMETERS_H_
`define PARAMETERS_H_

// `define col 16 // 16 bits instruction memory, data memory
// `define row_i 15 // instruction memory, instructions number, this number can be changed. Adding more instructions to verify your design is a good idea.
// `define row_d 8 // The number of data in data memory. We only use 8 data. Do not change this number. You can change the value of each data inside test.data file. Total number is fixed at 8. 
// `define filename "./test/50001111_50001212.o"
// `define simulation_time #160

localparam WIDTH = 32;
localparam REG_FILE_SIZE = 5;

`endif